// Maximum testing cycle
Bit#(32) maxCycle = 10000;

// Traffic Generator
typedef 10 InjectionRate; //Injection Rate: 0.XX
typedef 4 TrafficGeneratorSlotsCount;
